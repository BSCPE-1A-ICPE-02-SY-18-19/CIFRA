CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 39 210 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 1075 120 0 18 19
10 8 7 6 5 4 3 2 18 19
1 1 0 1 1 0 1 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3536 0 0
2
43530.4 0
0
2 +V
167 121 239 0 1 3
0 17
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4597 0 0
2
43530.4 0
0
9 2-In AND~
219 638 104 0 3 22
0 14 10 13
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3835 0 0
2
43530.4 0
0
9 2-In AND~
219 430 111 0 3 22
0 12 11 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3670 0 0
2
43530.4 0
0
7 Pulser~
4 66 414 0 10 12
0 20 21 15 22 0 0 5 5 4
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5616 0 0
2
43530.4 0
0
6 74112~
219 173 324 0 7 32
0 17 16 15 16 17 23 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9323 0 0
2
43530.4 0
0
6 74112~
219 343 323 0 7 32
0 17 12 15 12 17 24 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
317 0 0
2
43530.4 0
0
6 74112~
219 530 324 0 7 32
0 17 14 15 14 17 25 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3108 0 0
2
43530.4 0
0
6 74112~
219 700 323 0 7 32
0 17 13 15 13 17 26 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
4299 0 0
2
43530.4 0
0
6 74LS48
188 922 206 0 14 29
0 9 10 11 12 27 28 2 3 4
5 6 7 8 29
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
9672 0 0
2
43530.4 0
0
36
7 7 2 0 0 4224 0 11 2 0 0 3
954 170
1090 170
1090 156
8 6 3 0 0 4224 0 11 2 0 0 3
954 179
1084 179
1084 156
9 5 4 0 0 4224 0 11 2 0 0 3
954 188
1078 188
1078 156
10 4 5 0 0 4224 0 11 2 0 0 3
954 197
1072 197
1072 156
11 3 6 0 0 4224 0 11 2 0 0 3
954 206
1066 206
1066 156
12 2 7 0 0 4224 0 11 2 0 0 3
954 215
1060 215
1060 156
13 1 8 0 0 4224 0 11 2 0 0 3
954 224
1054 224
1054 156
7 1 9 0 0 4224 0 10 11 0 0 4
724 287
882 287
882 170
890 170
0 2 10 0 0 8320 0 0 11 14 0 3
592 288
592 179
890 179
0 3 11 0 0 8320 0 0 11 23 0 3
397 287
397 188
890 188
0 4 12 0 0 8320 0 0 11 25 0 3
211 288
211 197
890 197
0 4 13 0 0 8192 0 0 10 13 0 4
664 274
649 274
649 305
676 305
3 2 13 0 0 8320 0 4 10 0 0 4
659 104
664 104
664 287
676 287
7 2 10 0 0 0 0 9 4 0 0 4
554 288
606 288
606 113
614 113
0 1 14 0 0 8192 0 0 4 17 0 3
491 111
491 95
614 95
0 4 14 0 0 0 0 0 9 17 0 3
492 263
492 306
506 306
3 2 14 0 0 8320 0 5 9 0 0 4
451 111
492 111
492 288
506 288
3 0 15 0 0 8192 0 9 0 0 20 3
500 297
496 297
496 405
3 0 15 0 0 8192 0 8 0 0 20 3
313 296
309 296
309 405
0 3 15 0 0 4224 0 0 10 22 0 4
104 405
662 405
662 296
670 296
4 0 12 0 0 0 0 8 0 0 24 4
319 305
258 305
258 288
253 288
3 3 15 0 0 0 0 7 6 0 0 4
143 297
104 297
104 405
90 405
7 2 11 0 0 0 0 8 5 0 0 4
367 287
398 287
398 120
406 120
0 1 12 0 0 0 0 0 5 25 0 3
253 288
253 102
406 102
7 2 12 0 0 0 0 7 8 0 0 4
197 288
305 288
305 287
319 287
0 4 16 0 0 4096 0 0 7 27 0 4
39 288
135 288
135 306
149 306
1 2 16 0 0 8320 0 1 7 0 0 3
39 222
39 288
149 288
5 0 17 0 0 4096 0 10 0 0 36 2
700 335
700 351
5 0 17 0 0 0 0 9 0 0 36 2
530 336
530 351
5 0 17 0 0 0 0 8 0 0 36 2
343 335
343 351
5 0 17 0 0 0 0 7 0 0 36 2
173 336
173 351
0 1 17 0 0 0 0 0 10 36 0 2
700 248
700 260
1 0 17 0 0 0 0 9 0 0 36 2
530 261
530 248
0 1 17 0 0 0 0 0 8 36 0 2
343 248
343 260
0 1 17 0 0 0 0 0 7 36 0 4
174 248
174 253
173 253
173 261
1 0 17 0 0 4224 0 3 0 0 0 4
121 248
769 248
769 351
121 351
1
-16 0 0 0 700 0 0 0 0 3 2 1 66
11 Kristen ITC
0 0 0 28
327 472 588 507
338 480 576 503
28        Lord Devince S. Cifra
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
